library verilog;
use verilog.vl_types.all;
entity MAIN_vlg_vec_tst is
end MAIN_vlg_vec_tst;
