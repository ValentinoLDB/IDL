library verilog;
use verilog.vl_types.all;
entity validacionInicioFin_vlg_vec_tst is
end validacionInicioFin_vlg_vec_tst;
