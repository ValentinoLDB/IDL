library verilog;
use verilog.vl_types.all;
entity Prueba_vlg_vec_tst is
end Prueba_vlg_vec_tst;
