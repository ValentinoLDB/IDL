library verilog;
use verilog.vl_types.all;
entity CONTADOR_UPDOWN_vlg_vec_tst is
end CONTADOR_UPDOWN_vlg_vec_tst;
