library verilog;
use verilog.vl_types.all;
entity Sum_Res_vlg_vec_tst is
end Sum_Res_vlg_vec_tst;
