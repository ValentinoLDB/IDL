library verilog;
use verilog.vl_types.all;
entity validacionInicioFin_vlg_check_tst is
    port(
        error           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end validacionInicioFin_vlg_check_tst;
