library verilog;
use verilog.vl_types.all;
entity Sum_Res_vlg_sample_tst is
    port(
        A               : in     vl_logic_vector(11 downto 0);
        B               : in     vl_logic_vector(11 downto 0);
        Up_Down         : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Sum_Res_vlg_sample_tst;
