library verilog;
use verilog.vl_types.all;
entity Sumador1bit_vlg_vec_tst is
end Sumador1bit_vlg_vec_tst;
