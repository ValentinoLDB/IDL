library verilog;
use verilog.vl_types.all;
entity TPI_GRUPO03_vlg_vec_tst is
end TPI_GRUPO03_vlg_vec_tst;
