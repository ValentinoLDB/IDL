library verilog;
use verilog.vl_types.all;
entity MaquinaEstados_vlg_vec_tst is
end MaquinaEstados_vlg_vec_tst;
