library verilog;
use verilog.vl_types.all;
entity Contador_vlg_check_tst is
    port(
        Cont            : in     vl_logic_vector(11 downto 0);
        DATA            : in     vl_logic_vector(11 downto 0);
        sampler_rx      : in     vl_logic
    );
end Contador_vlg_check_tst;
