library verilog;
use verilog.vl_types.all;
entity Contador35_vlg_vec_tst is
end Contador35_vlg_vec_tst;
